module sound_artyx(
	input
);

endmodule