module tb_sound();
	

endmodule